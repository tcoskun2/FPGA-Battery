module topnet (
    input wire clk,
    input wire reset,
    
    output wire [31:0] predicted_soh
    
);
    //weights and biases concatenated in 32bit, Q16.16
    wire [32*4*64-1:0] weights1 = 'b11111111111111111101101000110000111111111111111110110101001100000000000000000000010110100001011011111111111111111010000101000110000000000000000000100111110110000000000000000000000100100001111111111111111111111110100011011111111111111111111111001010100011111111111111111111101101100110101100000000000000000010011000111101000000000000000000101111110100011111111111111111111110010001001011111111111111111001110101011101111111111111111110001100001111010000000000000000100001011000101000000000000000000111101001001001111111111111111111101111100010011111111111111111100011000110010111111111111111111111011010001001111111111111111111000111100110100000000000000000010010100011011011111111111111111011000000010101000000000000000000011100000000000000000000000000010010111101011000000000000000000111001010001110000000000000000000010001110110111111111111111111100110000111010100000000000000000111000010010010111111111111111111101000000000100000000000000000011000001100101111111111111111110110001100010101000000000000000001010000000110110000000000000000001111101110111100000000000000000001000010000110000000000000000000011010010110000000000000000000010101111001001011111111111111110111000101111110111111111111111110010111011111111111111111111111111101100100011000000000000000000101110000011100111111111111111110000111000110100000000000000000000011011100111011111111111111111010000101100111111111111111111111100110100101110000000000000000001011000100111000000000000000000110111111110100000000000000000001011111011101011111111111111111111110111110011000000000000000000111110001010011111111111111111111101110010000111111111111111111111110010000000100000000000000000000011100000100111111111111111101111100001110000000000000000000000111011001111100000000000000000101100001100100000000000000000001100110000001000000000000000000000010000010100100000000000000000101010100011001000000000000000000000111011111001111111111111111100001010010011111111111111111111101111100001010111111111111111110110011000010000000000000000000000110011000110011111111111111111101000100001010000000000000000001101000011111100000000000000000000010001110001000000000000000000101101101010100000000000000000000110000101001011111111111111111111111110110110000000000000000000101011001101001111111111111111111100111110010010000000000000000001111011001011000000000000000000111001010100001000000000000000001101111101011101111111111111111011101110111011111111111111111111001010101000011111111111111111111010101111000111111111111111111110101010011100100000000000000000100001011011101000000000000000000100101101000100000000000000000000001110111110100000000000000000100010001000110000000000000000001001111011000100000000000000000001101101111101011111111111111111110111011111000000000000000000010000000100000111111111111111111100111010101100100000000000000000000101101000010111111111111111101100010101100111111111111111111111110000101011111111111111111111111110000010111000000000000000000010111100100010000000000000000010111111000111111111111111111111011001001110111111111111111111110011111010000110000000000000000001110111100000111111111111111111111110100111101111111111111111111110000010101010000000000000000001101111111000111111111111111111010100000101010111111111111111110111111110011000000000000000000010100101011010000000000000000000011010001001101000000000000000001000010100101101111111111111111100111010101111011111111111111111001001001001010000000000000000000010110101001011111111111111111110100100011001111111111111111111001100110101100111111111111111111101000000000100000000000000000000001110101110000000000000000000110100110110000000000000000000010010100001000110000000000000000001000011010011011111111111111111010110000110111000000000000000000101100100110001111111111111111100100110111110011111111111111111111101100000100000000000000000000010011010110110000000000000000010000000001110011111111111111111101100100101000111111111111111111010011101000000000000000000000001000110110100011111111111111111110010010101110000000000000000001001010100000001111111111111111111011011101111100000000000000000001011011011011111111111111111110101100100110111111111111111111011010100011110100000000000000000100011101100111000000000000000010101101101000001111111111111111100101100010101111111111111111111000110000101000111111111111111110010111000010001111111111111111100000010011011000000000000000000101001100011011111111111111111110110100111011100000000000000000001010001011001111111111111111111001111101100110111111111111111110001011011011110000000000000000000000110000100100000000000000000110011011111101111111111111111111101010001011011111111111111111111101110111110111111111111111111010001000001101000000000000000000110010001000100000000000000000100010100101011011111111111111111011110100011001000000000000000010101101010100011111111111111111101100000000111011111111111111110111100111111011000000000000000010000011010000100000000000000000110010000101100011111111111111111110001100111100111111111111111110100101111000110000000000000000011101000100000100000000000000000011110101011110111111111111111111110011011011110000000000000000011101100001100111111111111111111101000011100101000000000000000001010001010101100000000000000000011010110101111011111111111111111111111000001100000000000000000001011111000010011111111111111111110110100011110111111111111111111000001101111010000000000000000001111101010000111111111111111111101010110011001111111111111111110010000001011111111111111111111111010110000100000000000000000000100011010101000000000000000000000000001100110110000000000000000000111011100110000000000000000000000101001000000111111111111111111100010001101011111111111111111111010000111111101111111111111111111001001000010011111111111111111110111111010001111111111111111110001100110110100000000000000000010100101000111000000000000000000110111010110010111111111111111110001101110000010000000000000000010000001001111000000000000000000000000000100001000000000000000001000001110011111111111111111111110011110110110000000000000000000101100101111001111111111111111110011110111000001111111111111111010001100000011100000000000000000100010010101101000000000000000001101001111001011111111111111111111101100001110100000000000000000000100110101010000000000000000001101101000101110000000000000000001111101111001000000000000000000000110011110001000000000000000001000001111110111111111111111111101001000101011111111111111111111100101010011100000000000000000000110000001010000000000000000000000010111101000000000000000000000011100101101100111111111111111111011100111010111111111111111111100010101011101100000000000000000010001010010000000000000000000001101100101111000000000000000000010111110100110000000000000000000101101101011111000000000000000010000001111111110000000000000000010100101010000111111111111111111001101110011000111111111111111110101100011010101111111111111111101000010001110011111111111111111011011000000110000000000000000001001010010001000000000000000000001010011011011100000000000000000110011010001101000000000000000000101111111000011111111111111111111101011100101111111111111111111111011010000000111111111111111111111111010111010000000000000000001010100010000111111111111111111001100001110001111111111111111110011000010000011111111111111111110001111111111011111111111111111101001101100111111111111111111111001100110001110000000000000000010011101110000000000000000000000100101100101111111111111111111110011000100000100000000000000000011110011100001111111111111111111010001001110010111111111111111111101111100010110000000000000000010101110011100111111111111111111110010111011111111111111111111111110010111101110000000000000000001110110001100011111111111111111011010100100001000000000000000000110110000110110000000000000000010001000011110100000000000000001101101100101111111111111111111111100011011101001111111111111111011100100100000000000000000000000110000011000101000000000000000000011101011110100000000000000000001111000111000011111111111111111011101101110101111111111111111111001000100010110000000000000000000001101000000011111111111111111101111011100110000000000000000001000000101100111111111111111111110010111101100000000000000000000010100010011000000000000000000000100011001001001111111111111111111111010011110111111111111111111001110010111001;
    wire [32*64-1:0] bias1 = 'b00000000000000000101110111100101000000000000000000110100100011101111111111111111011010010111001100000000000000000000100110111001111111111111111111011111111100101111111111111111100011001010001111111111111111111011001010001100000000000000000000101000111010001111111111111111111011111010110111111111111111111101001011110010000000000000000000000100100000000000000000000000010110111110101000000000000000000011000111110110111111111111111110110101100100101111111111111111100010111101011000000000000000000110100001101111111111111111111111101001010001111111111111111111100001110011110000000000000000000110000000010001000000000000000001010011000111010000000000000000000001100001101011111111111111111101001011010111000000000000000000100100000010101111111111111111100010100000101000000000000000000000010110101000000000000000000000101100110001100000000000000000010011010100011000000000000000000010001011000110111111111111111110001101011001011111111111111111110100011110100000000000000000000001011101000001111111111111111110011101001011101111111111111111111111101011111100000000000000000000101011110000111111111111111111011110011111100000000000000000000101101110101100000000000000000100111110100101111111111111111110011110000000001111111111111111111110110011010011111111111111111010000011100100000000000000000001110011001110111111111111111111110000001010101011111111111111111001001101111101111111111111111111100011001101001111111111111111101110110011010111111111111111111110111010011101000000000000000001111101100000010000000000000000000001000000011100000000000000000111100000101101000000000000000000011001100100001111111111111111110110100101100000000000000000000100100001101100000000000000000001011011110101101111111111111111011110100110000000000000000000000111010110000001111111111111111111101111001111111111111111111111110111010100010011111111111111111001010100101110000000000000000000110100011011000000000000000000011101100000111111111111111111111110001101010000111111111111111110110011110011100000000000000000001101110010011000000000000000000110111110010011;
    wire [32*32*64-1:0] weights2 = 'b1111111111111111111110001011010000000000000000000001010101100011111111111111111111100001000101100000000000000000000100101000001000000000000000000001011110001110111111111111111111101001011101110000000000000000000010100000011111111111111111111111011111100111000000000000000000100001010011000000000000000000000101010100010111111111111111111111100001010101000000000000000000011100000110111111111111111111111111100110001011111111111111111111110110001110111111111111111111001001110101011111111111111111111011010111000000000000000000000000100000110101000000000000000000000000010100000000000000000000000001001000010111111111111111111111110000010110111111111111111111101110110011110000000000000000000111100001111000000000000000000000100000000101000000000000000000011111101001101111111111111111111111011111110000000000000000000001101010000001000000000000000000000001110111110000000000000000000001000110011100000000000000000000000101000011000000000000000000000111010001110000000000000000000010110100110111111111111111111111100111100100111111111111111110100011011011110000000000000000000111111000111011111111111111111110111001001101000000000000000000010011000111101111111111111111101111010001111111111111111111111111100111010011111111111111111111101111010010101111111111111111111001000001111000000000000000000001111011111010111111111111111111100011110010001111111111111111110001010110011011111111111111111110011110110100000000000000000000101110001100101111111111111111111010010100001011111111111111111111001100110011111111111111111111100010110001001111111111111111111101111100011111111111111111111110101000110111000000000000000000011010010011001111111111111111111000100010110011111111111111111110001100111010111111111111111111100111001111110000000000000000000101110110100011111111111111111111111001100101111111111111111111111110001000111111111111111111111101100010000011111111111111111111000100000111000000000000000000011001010011110000000000000000000111010010010111111111111111111111110000100100111111111111111111110100110001101111111111111111111110010101010000000000000000000001110011001000111111111111111111111110011101011111111111111111111011000100111100000000000000000000110011111111111111111111111111111110001010001111111111111111111111011101000100000000000000000001100101001110111111111111111111101010011111001111111111111111111100001001010111111111111111111111111011110011000000000000000000010000001101000000000000000000000001110011010111111111111111111110010011010010111111111111111111100111010010111111111111111111111101100111000100000000000000000001011111010011111111111111111111100010110111011111111111111111111110100010101011111111111111111111100101111001000000000000000000000001000111000000000000000000000100001001100100000000000000000001101110010111000000000000000000011001001010111111111111111111111000110100111011111111111111111110011110000101111111111111111111100100100110100000000000000000000000101010001100000000000000000001010001011000000000000000000000001001101001101111111111111111111111100100001111111111111111111110001010000000000000000000000000000110000011110000000000000000000111010101111000000000000000000000110110011100000000000000000000000011111000101111111111111111111010101000100111111111111111111111011001100111111111111111111111111010010110101111111111111111111101110100111000000000000000000001110000110011000000000000000000000101011001010000000000000000000001100001111111111111111111111111111110111010000000000000000000000100011111000000000000000000000011001111010000000000000000000000011000000010111111111111111111111010111001100000000000000000000110101111101011111111111111111110010010011010000000000000000000001111000110111111111111111111111000000101000000000000000000000001011111111001111111111111111111110111111100010000000000000000000010101010110000000000000000000000000101001110111111111111111111110111010110100000000000000000000011101011011100000000000000000001110111001110111111111111111111110110111101111111111111111111111101100101011100000000000000000000001000100100000000000000000000000101100000000000000000000000000011010111111111111111111111111111111011100011111111111111111111110100111100011111111111111111111110010100001011111111111111111111001101011010111111111111111111001100101101011111111111111111111111101110011100000000000000000000001101100001000000000000000000101000000011010000000000000000001100010000010011111111111111111110110111010001111111111111111111001011110100010000000000000000000100010001111111111111111111111110101010011011111111111111111111100111101011111111111111111111111100001000011111111111111111111110010111110010111111111111111111101011010000011111111111111111111010101000110000000000000000000000011110001101000000000000000000011011000001111111111111111111110011101010111100000000000000000000110110001011000000000000000000110101001111010000000000000000000110110011101100000000000000000001011010000010111111111111111111100010000011110000000000000000000101010100011100000000000000000000111000100111111111111111111111101011000011010000000000000000000110000001101100000000000000000000011001011111000000000000000000011011010011110000000000000000000001101010101011111111111111111011010110101100000000000000000000000011110000010000000000000000000001010100000000000000000000000000100000100010111111111111111110110100001111000000000000000000001100100001010111111111111111111110110011011101111111111111111111110011111011100000000000000000000001000001100111111111111111111110001010101010111111111111111110101110110011110000000000000000000100100001001100000000000000000010000010110100111111111111111111111111011000100000000000000000000100011010011100000000000000000001000110010011000000000000000000011010011100000000000000000000000000011100000111111111111111111111001010011001000000000000000000001111001001000000000000000000000001011001011111111111111111111011111010011000000000000000000000010101011001011111111111111111111011010100101011111111111111111111010111111101111111111111111111101011101011110000000000000000000000101001110000000000000000000000010001101001000000000000000000101000000011111111111111111111111011111111000000000000000000000001111101001110111111111111111111110111110000110000000000000000000011001101001000000000000000000001011011110100111111111111111111110111101011101111111111111111111100110110000100000000000000000000000000110011111111111111111111100110101110100000000000000000000010100101100100000000000000000000111111000001111111111111111111101101110010001111111111111111111010110101011011111111111111111111110011000111000000000000000000010001110100000000000000000000000001101010010100000000000000000000000011111110000000000000000000000111101101011111111111111111111101000100000111111111111111111110100101101010111111111111111111101111010011110000000000000000000100011101101000000000000000000001011000101101111111111111111111011101000110000000000000000000000100110011001011111111111111111101111101001110000000000000000000011110100011110000000000000000000010010000010000000000000000000000010000100100111111111111111111101111001011001111111111111111110111010101000100000000000000000001011110111010111111111111111111100011111101011111111111111111111000100001100000000000000000000001100010010011000000000000000000001010111001010000000000000000000010101111001011111111111111111110010101100010111111111111111111100000100011010000000000000000000001101101111000000000000000000000110111110011000000000000000000010000011110000000000000000000000100001000001000000000000000000001010101000111000000000000000000001110010011110000000000000000000001011010010000000000000000000001101100101100000000000000000000010000100000000000000000000000000011011100001011111111111111111110110010011011000000000000000000001101100111000000000000000000000000101100111111111111111111111111010000101001000000000000000000000111110101101111111111111111110110111000000111111111111111111111000011101011111111111111111111110000111111001111111111111111111100101111001000000000000000000001000010100111111111111111111111111011010101010000000000000000000011000101110011111111111111111110011111011011111111111111111111101111100111011111111111111111111100011000111011111111111111111111111011101001111111111111111111110011101100111111111111111111111101010001111111111111111111111111101111001000111111111111111111111100010000101111111111111111111110011010101100000000000000000000011111010000111111111111111111100100000000011111111111111111111111000110100111111111111111111111011000000110111111111111111111011001100101010000000000000000000110101101010111111111111111111101010011100000000000000000000000010110101000100000000000000000000010000111010111111111111111111110110100010010000000000000000000000000110111001111111111111111111010111001011100000000000000000000001100101000111111111111111111100101000011011111111111111111110111101101111100000000000000000000010111010000000000000000000000011011111011000000000000000000000011011011111111111111111111111101111011111001111111111111111111110110100111011111111111111111111100010011110100000000000000000001101101010111000000000000000000010010111010111111111111111111111100101000100111111111111111111111010110111100000000000000000000000011000100100000000000000000000001111011011011111111111111111111110100111110000000000000000000001100110101000000000000000000000100111101101111111111111111111110110101011100111111111111111111100001010000010000000000000000000100111011010000000000000000000001011110101101111111111111111111111100011111001111111111111111111011100011001100000000000000000001110001000100000000000000000000011000110011100000000000000000000111000100100000000000000000000001001110011000111111111111111111100111111111011111111111111111111001110000101011111111111111111111011111010111000000000000000000000000011010010000000000000000000000110010000111111111111111111111111001011010111111111111111111101011111000101111111111111111111010110111110000000000000000000001110110001000111111111111111111101010001001111111111111111111111000000101101000000000000000000001000011011100000000000000000000001101010010011111111111111111111110010110000100000000000000000000111011111111000000000000000000000110011010010000000000000000000000101101000011111111111111111110010110000011111111111111111111011110000011010000000000000000000101110101001111111111111111111101100010000001111111111111111111100101110101110000000000000000000110001111011011111111111111111110110010011100111111111111111111111100010110110000000000000000000010010001001111111111111111111111000011100100111111111111111111100001100100001111111111111111111110110000011011111111111111111111000000100110000000000000000000011110111011000000000000000000000000101011000011111111111111111110011011000100111111111111111111101100000111110000000000000000000010110101110000000000000000000000010111010011111111111111111111100111100000100000000000000000000000100010111100000000000000000000011101011010000000000000000000010000111011010000000000000000000110010101110000000000000000000000010100010100000000000000000000000100010110101111111111111111111000100100010111111111111111111111101001101100111111111111111111110011000110011111111111111111111001001100001111111111111111111111000101101011000000000000000000001000000000111111111111111111111111011101101111111111111111111110000110000101000000000000000000010011011101010000000000000000000010001111100000000000000000000001001111111110000000000000000000011111110000100000000000000000000001010011111000000000000000000001100001100011111111111111111111111000111010011111111111111111111011011110001111111111111111111111010111010011000000000000000000011000100100110000000000000000000100010001001111111111111111111111111111010011000000000000000000000101011111111111111111111111111001111010000011111111111111111111110010000101000000000000000000001010111111001111111111111111111010000010101111111111111111111110011110101001000000000000000000000010111010000000000000000000000100011100010011111111111111111110010010100010111111111111111111111110110011100000000000000000000000101011100111111111111111111111001001010011000000000000000000011001000101011111111111111111111011000110111111111111111111111111001100010010000000000000000000011001000100001111111111111111111110001001101100000000000000000000110100011100000000000000000000011001011111001111111111111111111111000110111111111111111111111110001001000101111111111111111111111010100000011111111111111111111010110011001000000000000000000001000111000111000000000000000000000011110101101111111111111111111001111011011011111111111111111111110100100011000000000000000000000110001010011111111111111111111111111110011000000000000000000000010110101100000000000000000000001000000111011111111111111111111100000110101111111111111111111101011101000100111111111111111111100111001001001111111111111111111000111011111000000000000000000001110011010010000000000000000000001000101100001111111111111111111000011100110000000000000000000000110101101110000000000000000000000001111100100000000000000000000001101110001011111111111111111110010010000010111111111111111111110110100100111111111111111111110111101010001100000000000000000001011100100001000000000000000000010010000111101111111111111111111110011111000100000000000000000001111001110010000000000000000000001010000111010000000000000000000001010110101111111111111111111101011001110010111111111111111111100011001100011111111111111111111010110000111011111111111111111111000110011001000000000000000001001101111001000000000000000000000111000001010011111111111111111110011011010010111111111111111111111101110111000000000000000000010010111000100111111111111111111111011010100111111111111111111111101010101100111111111111111111111001110100101000000000000000000001010001011010000000000000000000010110111001000000000000000000001010000001111011111111111111111111011000000111000000000000000000000001000010010000000000000000000000111100110000000000000000000000010110001001000000000000000000100000111101001111111111111111111011011011111100000000000000000001011111001111111111111111111111111101100100000000000000000000000111001100010000000000000000000000010010000010000000000000000000011000011111110000000000000000000000011001011000000000000000000000001100100111000000000000000000001110001011101111111111111111111111100011010000000000000000000000111110001001000000000000000000010101100011011111111111111111101110010101011111111111111111111111110101110111111111111111111111110110101011100000000000000000000000001101101100000000000000000001000101011111000000000000000000010011110000110000000000000000000110001011010000000000000000000001101011010111111111111111111111101010001101111111111111111111111010111101110111111111111111111101111110011000000000000000000000011010110010000000000000000000000000100000011011111111111111111111001010000100000000000000000000101000000111110000000000000000000110000000100000000000000000000000010110001110000000000000000000000001100001100000000000000000000111110001011000000000000000000000001101100111111111111111111111100010100111110000000000000000000001101000000000000000000000000001101100111010000000000000000000001001000110011111111111111111111010000100111000000000000000000001100011000001000000000000000000001001011110010000000000000000000110010000010111111111111111111110101100001000111111111111111111110110001110101111111111111111111000011110011000000000000000000000010100011001000000000000000000010110011110000000000000000000000110101110010100000000000000000001010000101110111111111111111111110101000111110000000000000000001000110010110011111111111111111110101011101111000000000000000000110100110000010000000000000000000010111111001000000000000000000001010010001010000000000000000000001101100001111111111111111111111100110010011000000000000000000001000110111000000000000000000000000101000100101111111111111111111100001010000000000000000000000000111110000111111111111111111111110100101011101111111111111111110111111001101011111111111111111111111001001110000000000000000000000011000010001111111111111111111001011100111011111111111111111101111010111001111111111111111111111000001100100000000000000000001010010010011111111111111111111110011111010011000000000000000000100010011100011111111111111111111110111010011111111111111111111111001100001011000000000000000000011000101111010000000000000000000101111101011000000000000000000001000110000011111111111111111111110101001111111111111111111111111000011001111100000000000000000001100110111010111111111111111111111011000000010000000000000000000001000010011111111111111111111111111100000101000000000000000000010000001001111111111111111111111100101100000111111111111111111110011101000010111111111111111111100000111000000000000000000000000111110101000100000000000000000000000000010010111111111111111111101001011010111111111111111111111101001000101000000000000000000001100011001111111111111111111111111010011001010000000000000000000110011110101111111111111111111111111100000001111111111111111111111010111011100000000000000000000011010101101000000000000000000000010100101011000000000000000000000010001110110000000000000000000110001100110111111111111111111111010100101111000000000000000000010100110100100000000000000000000000100100011111111111111111111110101111011011111111111111111111100001111011001111111111111111111111111110100100000000000000000000000010001000111111111111111111111011101101111111111111111111111111100100101111111111111111111110011011010010000000000000000000001011101000101111111111111111111011111111001111111111111111111111000001010100111111111111111111100010101001101111111111111111111000101000011000000000000000000001000110011010000000000000000000011011111110111111111111111111110111101000000100000000000000000001110010110111000000000000000000011001111110010000000000000000000100100001010000000000000000000000110000100001000000000000000000011100101011110000000000000000000011101001100100000000000000000001101010100000111111111111111111101100101111011111111111111111111110000100110000000000000000000000111111110101000000000000000000000100011100110000000000000000000001011110110000000000000000000001000101000100111111111111111111111000000010011111111111111111111100011000001011111111111111111111000111110101111111111111111111110010101001110000000000000000000110111111100100000000000000000001110010101001000000000000000000001001010111101111111111111111111011101100101000000000000000000000000100101111111111111111111111100100011101101111111111111111111100100000110111111111111111111110100011111100000000000000000000000110011011101111111111111111110111111001110111111111111111111110011001111111000000000000000000001101010011000000000000000000000111111100110100000000000000000001101110101001000000000000000000001111101100001111111111111111111100011111111111111111111111111110010001000101000000000000000000011101101011001111111111111111111101011011111011111111111111111110000000010000111111111111111111111010101000011111111111111111111000111011001011111111111111111110001101011100000000000000000000001101110100110000000000000000000011001101111100000000000000000001000101110001000000000000000000001001100111101111111111111111111011010111000111111111111111111110100111011100111111111111111111110000111100101111111111111111111011011011010100000000000000000001111100000010000000000000000000011011101101100000000000000000000110111110111100000000000000000000110011000000111111111111111111111101010110100000000000000000000101100000001011111111111111111110110100110010000000000000000000001011111110111111111111111111111010011001010100000000000000000001000011001101000000000000000000010100000000011111111111111111111111010100110011111111111111111110000000100101111111111111111111110010010001100000000000000000000101011111100000000000000000000000110001101000111111111111111111100110011100111111111111111111111000011100101111111111111111111110010110011001000000000000000000000000000111101111111111111111111101110101001111111111111111111110110010101100000000000000000000010011111010010000000000000000000000110111100011111111111111111110000101111110000000000000000000000010000110111111111111111111111111010100001000000000000000000001111011110001000000000000000000010111000101011111111111111111111000100110011100000000000000000000010100011010000000000000000000001100011111111111111111111111111011110000010111111111111111111111001010100110111111111111111111100111110011010000000000000000000000110111100100000000000000000000110011010110111111111111111111101100110100001111111111111111111111101000111011111111111111111110001010101000111111111111111111100110011110011111111111111111111011000110101111111111111111111110010110110001000000000000000000011011011110101111111111111111111111000110101100000000000000000001101100100001111111111111111111110101111011001111111111111111111010110100010100000000000000000000000100000010000000000000000000001011110111000000000000000000000001010111001000000000000000000000101110111010111111111111111111111000100011111111111111111111111111111111010000000000000000000001001000010101111111111111111111111001010011110000000000000000000100001001010100000000000000000001011001010100111111111111111111100011000111001111111111111111111011000010001100000000000000000000010101111100111111111111111111101111110101110000000000000000000110101001010111111111111111111110001001001011000000000000000000001000001000001111111111111111111001100101101011111111111111111110111101010111000000000000000000011000010110001111111111111111111001110111010000000000000000000000101001011011000000000000000000001001101100000000000000000000000110001101110100000000000000000001010100001111000000000000000000001000001011111111111111111111111111101011011011111111111111111110101010010101000000000000000000010000110110000000000000000000000111011001111100000000000000000001111110011011000000000000000000010001111100011111111111111111111011011100010111111111111111111111110000011101111111111111111111110000010111101111111111111111111010110011000111111111111111111110110011110010000000000000000000001101001101011111111111111111111110110111110000000000000000000000001111101111111111111111111111111011101011100000000000000000000011011110110100000000000000000000000001000000000000000000000000011110110011101111111111111111111101111100110011111111111111111111111010001010000000000000000000001111011100010000000000000000000010100000000111111111111111111111110110001001000000000000000000011000101100000000000000000000000101001010001111111111111111111110000100001000000000000000000000010110001011000000000000000000000010111100100000000000000000000001101111101010000000000000000000001000101000001111111111111111111011110001110011111111111111111110010011101010111111111111111111110000011110111111111111111111111011011011011000000000000000000001001110000001000000000000000000000000001101110000000000000000000010100010011100000000000000000000001110000101111111111111111111011100101111101111111111111111111111111001111111111111111111111110011001110111000000000000000000010010010110100000000000000000000100001101001100000000000000000000111101110100000000000000000000001011110111101111111111111111111001110010011000000000000000000000101001011111111111111111111111110100111111110000000000000000000001111010110011111111111111111111010010111000111111111111111111101101011100101111111111111111111101101000100011111111111111111110001010011011000000000000000000100101011111100000000000000000000101011011111111111111111111111110001111011100000000000000000000010111111101100000000000000000000010001011110000000000000000000000010010100011000000000000000000000010100011000000000000000000000110101001100111111111111111111110101000110000000000000000000000010111111110101111111111111111111101001111111011111111111111111111111001111101111111111111111111110101001110110000000000000000000010110001110111111111111111111101011100001011111111111111111111100110111100000000000000000000000001000001010011111111111111111110111001000010111111111111111110100110000101110000000000000000000100010010001100000000000000000000011100010000111111111111111111110010011001101111111111111111111110110110101000000000000000000000001111001100111111111111111111000100110100101111111111111111110111001101011100000000000000000000000010001010111111111111111111110000011000010000000000000000000101000000011000000000000000000000010010010101000000000000000000010011111000000000000000000000000001000000011000000000000000000000010111101011111111111111111111111000010011101111111111111111111101100110101111111111111111111100111111110010000000000000000000001100010000010000000000000000000001000011110100000000000000000001011000000010000000000000000000010011001000000000000000000000000100001011100111111111111111111111000111011100000000000000000000100100111010001111111111111111111110100110111000000000000000000000100110011001111111111111111111101101111000011111111111111111111011110111000000000000000000000001100011101010111111111111111111101110110000001111111111111111111001110101100111111111111111111110101110010110000000000000000000001111101011100000000000000000000000110010111111111111111111111110000000110011000000000000000000011011011001011111111111111111111001011100100000000000000000000001000111111010111111111111111111101110101010000000000000000000000100100000000100000000000000000001110110000100111111111111111111111101110010011111111111111111111000011100110100000000000000000000010010000110111111111111111111101011001001011111111111111111111111011001001011111111111111111110110011001111111111111111111111111010001100000000000000000000000000111110110000000000000000000001001001100110111111111111111111100001011010110000000000000000000111101011010111111111111111111111111110000011111111111111111111111111000110000000000000000000000101010110101000000000000000000000001000011101000000000000000000011001010101001111111111111111111101001110001000000000000000000000101111010100111111111111111111111100111010101111111111111111111101110011100011111111111111111110100000000101000000000000000000001000111110101111111111111111111101100100000000000000000000000000011011111101111111111111111111100100011001000000000000000000000010111000100111111111111111111110101000101101000000000000000000011000110010011111111111111111111101010111100011111111111111111111100001010010111111111111111111111010011000111111111111111111111111001101101011111111111111111110010001000110111111111111111111101010011011011111111111111111111001100011011111111111111111111110111010111000000000000000000000000001110000100000000000000000000111001100010100000000000000000001011011001000111111111111111111111101101001111111111111111111111011001010100011111111111111111110111110011001111111111111111111100111111001001111111111111111111000001011110100000000000000000001001100010011111111111111111111100011001111100000000000000000000010101010110111111111111111111111111000011010000000000000000000000111000010011111111111111111111101111100011100000000000000000000101110010111000000000000000000010110100111111111111111111111111111111011011011111111111111111101111011101011000000000000000000010001101001101111111111111111111000110111101100000000000000000000100100001100000000000000000000011010011001100000000000000000000111000100111100000000000000000000111000110001000000000000000000010101001101111111111111111111111110011110101111111111111111111110000110110111111111111111111111110000110001001111111111111111111000110100110000000000000000000000100101101010111111111111111111101111010010011111111111111111111111101101011011111111111111111110111001000010000000000000000000001010110011101111111111111111111111110010100111111111111111111111101001010001111111111111111111101011110110001111111111111111111001110111001100000000000000000001111111010101111111111111111111111100010010001111111111111111111000001110101011111111111111111110100011101101111111111111111111101100000011000000000000000000000001110000111100000000000000000001111010011010000000000000000000001001011001011111111111111111111001111101101111111111111111111110011001000001000000000000000000001010101000110000000000000000000110110011001011111111111111111110010011100010000000000000000000010100111010101111111111111111111101101000000111111111111111111110001100110010000000000000000000011010000001101111111111111111111111110100110011111111111111111110111101001001000000000000000000000110000000011111111111111111111011001000011100000000000000000000010000001011111111111111111111111011110000111111111111111111111100100110100111111111111111111111010011001110111111111111111111110100010110000000000000000000000001111111001000000000000000000000001111001111111111111111111111101011010101110000000000000000000001010110010011111111111111111110101100110111000000000000000000001100001101000000000000000000000101001101001000000000000000000001010011100000111111111111111111110001011010001111111111111111111000101101000111111111111111111110101010111111111111111111111111100110101101000000000000000000000110001100000011111111111111111110000010111111000000000000000000000100010101011111111111111111111010001001011011111111111111111111010011000111000000000000000000100100010100101111111111111111111011101110100100000000000000000001010111110001111111111111111111110010101111011111111111111111111100110101000000000000000000000000000110110100000000000000000000011001110000011111111111111111110101100110111000000000000000000000110001111001111111111111111111101111101001000000000000000000000000100001110111111111111111111110110101001000000000000000000000010111010011000000000000000000000111110100011011111111111111111111011101001000111111111111111111010011110101000000000000000000001001000100101100000000000000000001100010100011111111111111111111110110111000101111111111111111111011110110101000000000000000000001100001111011111111111111111111100110001111110000000000000000000110010101001100000000000000000001110001101011000000000000000000001010101011001111111111111111110110010101000000000000000000000000100010110001000000000000000000001100011100111111111111111111111011100110000000000000000000000101000000000101111111111111111111101110010100100000000000000000000010011000000111111111111111111111010101011101000000000000000000101011011000011111111111111111110010100110101111111111111111111110110100111011000000000000000000011100100010010000000000000000000000101010000011111111111111111110001101010100000000000000000000110101111101001111111111111111111000101101000100000000000000000000001111011111111111111111111111101110001011001111111111111111111110000110001100000000000000000001101011011110000000000000000000011010111011111111111111111111111011011001011011111111111111111111000100111101111111111111111111110101001000011111111111111111111011100010001000000000000000000010100101001001000000000000000000001000101000111111111111111111111100100000110000000000000000000000110010010100111111111111111111100010011011001111111111111111111010001110011000000000000000000000011100001010111111111111111111000111111010011111111111111111111000001100001000000000000000000000001011111101111111111111111111100101010011000000000000000000000110101110111100000000000000000000011101101100000000000000000000001010001010011111111111111111110100010000001011111111111111111111101000110011111111111111111111110101001101100000000000000000000101100110010111111111111111111111111011111110000000000000000000001110010011100000000000000000000001001110111111111111111111111110111100110000111111111111111111110010010011011111111111111111111100001110001100000000000000000000110011011110111111111111111111110101011011001111111111111111111000111000001100000000000000000000101000100111000000000000000000100001100010110000000000000000001100101101010111111111111111111111100110101000000000000000000000010010011101010000000000000000000001001111110011111111111111111110100110101101000000000000000000001011011000100000000000000000000111000101110111111111111111111110101111111101000000000000000000011000011000000000000000000000000000111111001000000000000000000001000101111101111111111111111111111111001010110000000000000000000010001110101100000000000000000001001010110100111111111111111111000101100010111111111111111111111101000001101100000000000000000001100010010110000000000000000000010011111111101111111111111111101101001000100100000000000000000010011111111101000000000000000000001100101001111111111111111111111101010110011000000000000000000000001101000101000000000000000000000100101000011111111111111111100101010101101111111111111111111111110011011100000000000000000000110001011101110000000000000000000110011101001100000000000000000001000001010110111111111111111111011111110100011111111111111111110111001110001000000000000000000000110101101010111111111111111111100110001010000000000000000000000010100001101000000000000000000001101010110001111111111111111111011000111110001111111111111111111000110010000100000000000000000000000011100010111111111111111111110110110000110000000000000000000100010100001100000000000000000001101101000010000000000000000000000101111001100000000000000000010100101011110000000000000000000000001010011011111111111111111111111000101000011111111111111111110110101011000011111111111111111110000000011100000000000000000000000111101100111111111111111111111100101101111000000000000000000001101110111010111111111111111111111001010101010000000000000000000000110110010100000000000000000000000110111110111111111111111111101101100000101111111111111111111111110100100011111111111111111111011100111011111111111111111111111010110111000000000000000000000000010111110111111111111111111111000000000001111111111111111111110011010001011111111111111111111110001000011000000000000000000001011011111010111111111111111111111100111100111111111111111111111001011110001111111111111111111110000111010101111111111111111111100010000010001111111111111111111001000110101011111111111111111110111100011001000000000000000000001100110110010000000000000000000011010010010100000000000000000000110111110011111111111111111111111011110100010000000000000000000001010101110011111111111111111111011110000010000000000000000000001011010101110000000000000000000011111110111000000000000000000001011100110110000000000000000000010110000100100000000000000000000110011010100011111111111111111111100001100111111111111111111111101010010010110000000000000000000011010011010000000000000000000001111110010110111111111111111111110010011010010000000000000000000100101110101011111111111111111110101010000010111111111111111111110101011110100000000000000000000100100001101111111111111111111110101001111110111111111111111111101100011000010000000000000000000011111100111100000000000000000001101100101000111111111111111111100111010000000000000000000000000111110010000100000000000000000001100011000111000000000000000000000011000111011111111111111111111001100011010011111111111111111111010110001101000000000000000000000011101011000000000000000000000011111100100000000000000000000001110000110100111111111111111111101100001000010000000000000000000111111101001111111111111111111110101000011001111111111111111111100100110001100000000000000000000101100010110011111111111111111110101100001100000000000000000000010000101011010000000000000000000000010010011111111111111111111110011001010010111111111111111111110011101011001111111111111111111110111100000000000000000000000000000110111000111111111111111111100110100010011111111111111111111101011100011100000000000000000000001010001011111111111111111111111101101000000000000000000000000010000011000011111111111111111110111010100001000000000000000000011000111111110000000000000000000001001010100000000000000000000000001010001110000000000000000000011010111101111111111111111111111001110000001111111111111111111111100100110000000000000000000000001001110000010000000000000000000001101111001000000000000000000000011010110010000000000000000000000101000110011111111111111111111110011000011111111111111111111111001000101000111111111111111111110101111010011111111111111111111101111110101100000000000000000001111010100110111111111111111111100011001001110000000000000000000100111010001100000000000000000000011111101010000000000000000000000001100011111111111111111111111010011011000011111111111111111110001111000000111111111111111111111111011010000000000000000000000100100000000111111111111111111110111010011001111111111111111111101011001100001111111111111111110111111010111100000000000000000001011111010101111111111111111111111001110000101111111111111111111101000010101100000000000000000001000111111111111111111111111111101000110110010000000000000000000011110101001100000000000000000001000110100111111111111111111111101011000011011111111111111111111101110111001111111111111111111111100000110101111111111111111111100000110000000000000000000000000001101101111100000000000000000000000000100011111111111111111111111010000000001111111111111111111101111000011111111111111111111111011011101101111111111111111111101000100000110000000000000000000001011101001000000000000000000000000011001111111111111111111111110111010100001111111111111111111001010101110011111111111111111111111000000110111111111111111111101100101101010000000000000000000001110111101100000000000000000000111010001110000000000000000000011110000011001111111111111111111110111100101100000000000000000000001011011100111111111111111111110010011001111111111111111111111010100000101111111111111111111111010101010100111111111111111111110011101010001111111111111111111110100101110111111111111111111111101010100000111111111111111111111010100101110000000000000000000110110110001111111111111111111111000011111001111111111111111111110011100101001111111111111111111001001110111000000000000000000000011000100100111111111111111111101000101001100000000000000000000010001011101000000000000000000000010011001001000000000000000000001010001100001111111111111111111000100101101011111111111111111110110010110100111111111111111111101100000001101111111111111111111101100110100100000000000000000000100011110011111111111111111111111010000110001111111111111111111010101010111011111111111111111111011101000110000000000000000000011011110011110000000000000000000000110011011011111111111111111111000000010111000000000000000000011011101100010000000000000000000000001011001100000000000000000001101010011100000000000000000000010011110001001111111111111111111101111000001011111111111111111111100101010110111111111111111111110100000111110000000000000000000101111111110011111111111111111111000101010011000000000000000000010000110100000000000000000000000111100111100100000000000000000001001001000110111111111111111111101111001110000000000000000000000011110110001011111111111111111111001100110101000000000000000000011001101111000000000000000000000110001101111000000000000000000000111011111101111111111111111111110100001100010000000000000000000000101011110111111111111111111111111001000101000000000000000000000100000000001111111111111111111100101000111111111111111111111110110001001101111111111111111111110100111101011111111111111111111000110001111000000000000000000000001101011010111111111111111111110000101011111111111111111111111011111110001011111111111111111111011100110011000000000000000000010011000010111111111111111111111001111010000100000000000000000000100111010001000000000000000000010100011001111111111111111111111011100110001000000000000000000001001011001111000000000000000000011111100101000000000000000000000001110110000000000000000000000001111111011111000000000000000000000000000101100000000000000000000010110111111111111111111111111110110010001011000000000000000000010100111101100000000000000000000100001110101000000000000000000000001010100101000000000000000000101100111001010000000000000000000101100100100011111111111111111110111011011011000000000000000000000011011001000000000000000000000010110110100111111111111111111101111101110001111111111111111111111001100110001111111111111111111101001101111100000000000000000000000101111010000000000000000000000011010100100000000000000000000011110110100100000000000000000001101110110110111111111111111111110010100001101111111111111111110111111001100111111111111111111111100010011001111111111111111111101010111011010000000000000000000001100001100111111111111111111110011000010101000000000000000000010110001101101111111111111111111000100010111011111111111111111111001011011110000000000000000000011000101111011111111111111111111010100101111111111111111111111111011110001110000000000000000000011101000101001111111111111111100011000111000011111111111111111110110011110111000000000000000000000100110100100000000000000000000000010101101111111111111111111001011101001111000000000000000000010011100110000000000000000000000000111100111000000000000000000000110100001010000000000000000000001000100101011111111111111111111000000001001111111111111111111010011111110011111111111111111111101100100110010000000000000000001111001101001111111111111111111110010001101100111111111111111111111111100101010000000000000000000011111001101100000000000000000001100000000000111111111111111111111101110010111111111111111111111001010001010011111111111111111110001010100000000000000000000000011000000001001111111111111111111000011011000100000000000000000000110010001001000000000000000000001010110100111111111111111111111101010000101111111111111111111110100110100100000000000000000000001110101010101111111111111111111110101101000100000000000000000101001110000011111111111111111111111101110110010000000000000000000111111111001011111111111111111110111010001011000000000000000000000111100110010000000000000000000001110010010000000000000000000001000101101110111111111111111111011100010011000000000000000000000111100100001111111111111111111101110100010100000000000000000000011111110100000000000000000000000110000110001000000000000000000000010000000011000000000000000000010100000110001111111111111111111011001100101111111111111111111111110011010100000000000000000000010101011110101111111111111111111101110110100111111111111111111101011101110000111111111111111111110110100110110000000000000000000010100100101000000000000000000000001101011100000000000000000000001101111101000000000000000000000100110001111100000000000000000001010011001110000000000000000000000000110000000000000000000000000100100001101011111111111111111111010011101100111111111111111111100101111001110000000000000000000100010010000011111111111111111111100101101010000000000000000000010101100011001111111111111111111100000001000111111111111111111111011010101000000000000000000000010001001011100000000000000000000010010100011011111111111111111101100101101010111111111111111111101111011010010000000000000000000001100100010100000000000000000001011111110101111111111111111110110000010101100000000000000000000111010000101000000000000000000000111000100101111111111111111111100110111011010000000000000000000110101000101011111111111111111110001110111111111111111111111110110000011110011111111111111111111110101100110000000000000000000001100100110101000000000000000000000001001000110000000000000000000110000100100111111111111111111110000011011010000000000000000000001110010010010000000000000000000001011010010111111111111111111111011011010100000000000000000000010110001010111111111111111111111110100001000111111111111111111110001111100110111111111111111111101111101010101111111111111111110111100100110000000000000000000001000001011011111111111111111111110011110101101111111111111111111001111111101100000000000000000000100011100110000000000000000000001101101100011111111111111111111101010101110111111111111111111111110101000001111111111111111111110011100111100000000000000000000000100001001111111111111111111101110001110011000000000000000000001110111110000000000000000000000101100100011000000000000000000001001010011010000000000000000000010001110001010000000000000000000001100000101100000000000000000000101101011110111111111111111111111111011100101111111111111111110111000001100011111111111111111110010101110100000000000000000000100001111100001111111111111111111001001010100100000000000000000000010111001100111111111111111111111100001001111111111111111111111100000101010011111111111111111111001110001110111111111111111111110100110100110000000000000000000010011010110000000000000000000000001010001000000000000000000000001011111010100000000000000000000010010111001100000000000000000001001100111010000000000000000000001100011001010000000000000000000011000000101111111111111111111111001111001111111111111111111111100000001110011111111111111111111101001011100000000000000000000000110110010101000000000000000000000111011000011111111111111111111000100110001011111111111111111110011101010101000000000000000001001011010101110000000000000000000011100110001011111111111111111111011011010101111111111111111111011110000111110000000000000000010010001000011111111111111111111101111110111001000000000000000000001011010110000000000000000000000110000011110111111111111111111110110011100010111111111111111111100000111011000000000000000000000101110010111011111111111111111110011000110011111111111111111111110111100100100000000000000000000100010011000000000000000000000001011101101101000000000000000000000100101111000000000000000000000101000110000111111111111111111111101100101000111111111111111111100001011100000000000000000000000100000000010111111111111111111110110000000101000000000000000000011010110011110000000000000000000111111001000011111111111111111111101101101010111111111111111111100100101011101111111111111111111010001101111111111111111111111111011000011111000000000000000000001111110001001111111111111111101100101110010011111111111111111111010010010001111111111111111111101001101001011111111111111111111001101001001100000000000000000001100001111011111111111111111111110001001010010000000000000000000000101001110011111111111111111111011100101110000000000000000000000110000000001111111111111111111110101100000000000000000000000000010100011011000000000000000000100110111111101111111111111111111010110011101100000000000000000000010100111111111111111111111111111001110000001111111111111111110111111110110100000000000000000001100001111110111111111111111111110010110001111111111111111111111011000011100100000000000000000000000100101001000000000000000000000010000000001111111111111111111111010010110000000000000000000001000000001101111111111111111111100001011111101111111111111111111010110100000111111111111111111111111011100010111111111111111111101001101001011111111111111111111100000111001011111111111111111111111011101011000000000000000000010100111010001111111111111111111011111001010111111111111111111111011000011100000000000000000000101010001100010000000000000000000000101101111100000000000000000001010110011101000000000000000000010101010100011111111111111111101100101111111011111111111111111111010001111001111111111111111111011010000000000000000000000000000011101001111111111111111111111001101111100011000000000000000000101110100110100000000000000000001010101011011000000000000000000000000010000101111111111111111111110010101100001111111111111111111111111101101011111111111111111000100110010010111111111111111111110000001111000000000000000000001101001001000011111111111111111111001110111111111111111111111111100010010001110000000000000000000000000110100100000000000000000001101011001111000000000000000000001001000001100000000000000000000011110110001100000000000000000001010111001011111111111111111111110100011101011111111111111111111011010101100100000000000000000000101101000111111111111111111111101110100010100000000000000000000010111101101100000000000000000000111010010000000000000000000000011001111000001111111111111111111100001101011100000000000000000010111101101010000000000000000000100110000111010000000000000000000001000001110011111111111111111111100011011011111111111111111111111000010001011111111111111111111111110000111011111111111111111111110101101110000000000000000000010010100001001111111111111111111000111011111111111111111111111110111100011100111111111111111111110010001001110000000000000000000101100111111000000000000000000000011001000010111111111111111111111000100110010000000000000000000101001100001100000000000000000000111101100000000000000000000000000000000000100000000000000000000101010100011011111111111111111111111010001000000000000000000000000010100111010000000000000000000001000101100100000000000000000001111110100010000000000000000000011000011000011111111111111111111011111110011011111111111111111110010000001101000000000000000000001010111101100000000000000000000001011000000100000000000000000000110101110010000000000000000000001000111101101111111111111111111010001111010111111111111111111110111101100001111111111111111111111010011011100000000000000000000000001100100011111111111111111111111010101111000000000000000000001100100101111111111111111111111001100110101011111111111111111010111010000010111111111111111111110000011010111111111111111111111111010100001100000000000000000010000011110101111111111111111110110000001011001111111111111111111110000010011100000000000000000001011001110101111111111111111111111010000010001111111111111111111001110001010011111111111111111110000011111110111111111111111110111011101001001111111111111111111111001100001111111111111111111111011100011000000000000000000000010100011111001111111111111111111001101000001100000000000000000000010011011011000000000000000000001000011100001111111111111111111100111111010011111111111111111111111011011000000000000000000000010001110101010000000000000000000110011000111100000000000000000000101011100110000000000000000000000010011011001111111111111111111111100001001000000000000000000001001110101011000000000000000000000011011010011111111111111111111001110100001011111111111111111111101100011111000000000000000000110111001111111111111111111111111101001001011000000000000000000001101110101110111111111111111111100001100100111111111111111111111000001111110011111111111111111111101110100011111111111111111111110000100001010000000000000000000110110101101000000000000000000001011011010110111111111111111111111010111010101111111111111111111111001011000011111111111111111111000010001011000000000000000000001000000010011111111111111111111100011010000111111111111111111111010011110111111111111111111111111110001100001111111111111111111110011001010011111111111111111111011010110010000000000000000000001100001111111111111111111111111000101100001111111111111111111110010001111001000000000000000000000011101001000000000000000000000000100010111111111111111111111110011010110110111111111111111111100000110111010000000000000000000010100110100000000000000000000001100011001110111111111111111111110100001000101111111111111111111110111101011000000000000000000000111100100011000000000000000000001001110101011111111111111111111100001001100100000000000000000000010111000000000000000000000000011011110000111111111111111111111101001101101011111111111111111111010010100000111111111111111111110100000010100000000000000000000000000110000000000000000000000000000100000000111111111111111111101100010010110000000000000000000011110011100011111111111111111110011101011100111111111111111111100000001001001111111111111111111101100011101111111111111111111111100100100110000000000000000000011001010011001111111111111111111010010001110011111111111111111110001000011111111111111111111111100000011100100000000000000000000011111110100100000000000000000001001010101000111111111111111111111101001101101111111111111111111011011101000000000000000000000001001111101111111111111111111111110010111000100000000000000000000000010101011000000000000000000001100110110011000000000000000000000101001101000000000000000000000010011000101100000000000000000000111000011011111111111111111111111010010100011111111111111111111010010100111000000000000000000000001011011101000000000000000000011100001010110000000000000000000011110000000000000000000000000000000011100001111111111111111111101101001011001111111111111111111001011110100100000000000000000000011000100111000000000000000000001000001100110000000000000000000101010111001011111111111111111110111110101100000000000000000000011101110000110000000000000000000110101010111011111111111111111111000101111000111111111111111111111100011001111111111111111111111101101101100100000000000000000000000000000000111111111111111111100110010001111111111111111111111000010011111011111111111111111110100000001111111111111111111111111010001110011111111111111111111111110011100000000000000000000001100100110010111111111111111111100011100100111111111111111111111010110100011000000000000000000001111010010000000000000000000000000001100111011111111111111111111010001010010100000000000000000001011111011100111111111111111111100111101010011111111111111111111111010101100100000000000000000000000010011000000000000000000000000111011001111111111111111111111000110000100000000000000000000001111001010010111111111111111111111101011110100000000000000000000011010100100111111111111111111110101111001100000000000000000000001001100011001111111111111111111011011010110100000000000000000001111000110010111111111111111111101101010001101111111111111111111010101010110100000000000000000001110010011100111111111111111111111001110011000000000000000000000111010010101111111111111111111110001100011001111111111111111111110011100000110000000000000000000010101000110100000000000000000000010100001111000000000000000000011011001111111111111111111111111100001011101000000000000000000000011011100001000000000000000000001111011001101111111111111111111000000100001000000000000000000001100001110011111111111111111111100010101111110000000000000000000010100111011111111111111111111110100111101110000000000000000000011001101001011111111111111111111111110100111000000000000000000000000001101011111111111111111111101001011101100000000000000000000001100100011011111111111111111111100001000001000000000000000000011011010001011111111111111111111011001000101011111111111111111111011101100010111111111111111111111101110110001111111111111111111110010000100111111111111111111111101111010101111111111111111111101001101001100000000000000000000010010100101000000000000000000000000100101110111111111111111111110010101101111111111111111111111011101110101011111111111111111111001100010111000000000000000000011010011100011111111111111111111101011010110011111111111111111110011001111110111111111111111111101101001100111111111111111111111000011000001000000000000000000000101011001111111111111111111111100010101110101111111111111111111001101110000100000000000000000000000010100001000000000000000000001001001100101111111111111111110111110100000000000000000000000000100010000001000000000000000000001100000111001111111111111111111111111110010100000000000000000001100000110111111111111111111111101100010010101111111111111111111010010110010000000000000000000000100100010111000000000000000000010011100111000000000000000000000101000110011111111111111111111110000111010101000000000000000000011100111001100000000000000000000110011010100000000000000000000001011010111001000000000000000000001010010001111111111111111111111101110110110111111111111111111110001000111010000000000000000000000001111100101111111111111111110111100111110100000000000000000001100101111000111111111111111111011011011111100000000000000000000101110011011000000000000000000010011001110011000000000000000000010101000011010000000000000000000010101100011000000000000000000000000001111011111111111111111111000101000101011111111111111111111011111110011000000000000000000001010110110100111111111111111111110100100100001111111111111111111001001001111011111111111111111110001100100010111111111111111111111101101010000000000000000000000101101000100111111111111111111110100000101011000000000000000000011011101011111111111111111111111001111110011011111111111111111111101010000110000000000000000000000010111001110000000000000000000101010110111100000000000000000000110100001010111111111111111111110111010110001111111111111111111001000111000000000000000000000000001110010000000000000000000000011100100110000000000000000000000101111000000100000000000000000000110011100001111111111111111111111000001010100000000000000000000011110010011000000000000000000001110100010111111111111111111111101000111110000000000000000000000101011100110000000000000000000000100101011000111111111111111111101111010110110000000000000000000010111001001100000000000000000001010001100000000000000000000000001010100011100000000000000000000001010101011100000000000000000000010111001111111111111111111111101110111101010000000000000000000010001100000111111111111111111111001101101111000000000000000000001001001101001111111111111111111011110011011011111111111111111111011110001010000000000000000000011010101010111111111111111111111110001111011100000000000000000000100101011010111111111111111111111100111100101111111111111111111100011011000011111111111111111111011010011100000000000000000000001001110101001111111111111111111110010101010011111111111111111110011101111010111111111111111111111100001101011111111111111111111001001110011111111111111111111110000110111100111111111111111111110100000100000000000000000000000111100100000111111111111111111110000110000101000000000000000000001101111101011111111111111111111101011000110111111111111111111110010111101100111111111111111111111010000110000000000000000000000001010001000000000000000000000000100111101010111111111111111111111000101001000000000000000000000011000101001011111111111111111110110001101010000000000000000000001011110000010000000000000000000100111110000111111111111111111111001111010011000000000000000000010010001100101111111111111111111111010000101000000000000000000000011101010111000000000000000000000001010001011111111111111111111000011000111100000000000000000000010111011111111111111111111111111110010001001111111111111111111010011100010100000000000000000000101000111001111111111111111111110101000001011111111111111111111101010110001100000000000000000000111001110010000000000000000000011001101001100000000000000000000010000111100011111111111111111110000111011001111111111111111111100110111101100000000000000000000100111101111100000000000000000001001101100011000000000000000000000010001001110000000000000000000101011000100011111111111111111111010011000110111111111111111111100101011110001111111111111111111001001010111111111111111111111111000110110001000000000000000000001100111010111111111111111111111101101101011000000000000000000000101110110000000000000000000000010111001101100000000000000000001000010100000111111111111111111110001111001101000000000000000000011100000101001111111111111111111011100101011011111111111111111111111001010000111111111111111111111100010101101111111111111111000101111001111100000000000000000000010100001110000000000000000000001010101001101111111111111111111100000101101000000000000000000000011101101011111111111111111111100011111111110000000000000000000001100011101100000000000000000001011000110110000000000000000000001100010110111111111111111111111000110111111100000000000000000000010001100001111111111111111111111100100011111111111111111111111001110011110100000000000000000001001111000011000000000000000000011000010110010000000000000000000011111001010011111111111111111110000010001000000000000000000000010011101011111111111111111111011000100001010100000000000000000001011100001110111111111111111111100000100110101111111111111111111011100001100111111111111111110110011111100011000000000000000000101100111100010000000000000000001010100011110011111111111111111111100001000101000000000000000000011111111000011111111111111111111111111111000111111111111111111001101001110101111111111111111111111011111001011111111111111111111111110110000000000000000000000001001000110011000000000000000000000001111101001111111111111111111010100101100000000000000000000001101100011010000000000000000000000100111000101111111111111111111110000011010000000000000000000001000001001001111111111111111111111111100010101111111111111111110101110100010011111111111111111111100111010111000000000000000000000110001010100000000000000000001000101000101000000000000000000001011111010100111111111111111111110000001101110000000000000000000101000100010000000000000000000101000001010101111111111111111110011110001100101111111111111111111011001101010000000000000000000000110000010111000000000000000000001100000111001111111111111111111100100001010100000000000000000000010111100000111111111111111111101100100101111111111111111111111011100100011000000000000000000000111011110100111111111111111111111101100011110000000000000000000010100110001011111111111111111111011111110101000000000000000000011101000110101111111111111111111011000011010100000000000000000000101101000011000000000000000000000110100101011111111111111111111011111011101100000000000000000001011111101010000000000000000000000101111101001111111111111111111100011010101011111111111111111111011100100111000000000000000000010010010111001111111111111111111110000111011000000000000000000000010110101111000000000000000000101100000111000000000000000000000111000011000011111111111111111110010010001000000000000000000000011100110101001111111111111111111100001100110100000000000000000001011001001010111111111111111111101100111111000000000000000000000011001011001011111111111111111111101100001010000000000000000000001001000010111111111111111111111011100110100111111111111111110111100010001101000000000000000000010101110101000000000000000000000100000100000000000000000000000001100011000100111111111111111110110101110111110000000000000000010100101010011100000000000000000001011010101010000000000000000000011111111100010000000000000000000010011100010100000000000000000000010101111000111111111111111110000111000110100000000000000000000011010110011000000000000000000011101111010110000000000000000000000101110001010000000000000000000001110110110111111111111111111110011011010010000000000000000000001101100000110000000000000000000110111101010011111111111111111111000111110010000000000000000000001111011011011111111111111111111010110010110111111111111111111011010100111110000000000000000000100001011000001111111111111111111001000000111011111111111111111111101001100111000000000000000000000101001001100000000000000000001000110010110111111111111111111110101001001010000000000000000001011010110101111111111111111111111010001001100111111111111111111111011010001100111111111111111111100110010010010000000000000000000000001010010100000000000000000000001101111001111111111111111111100110000001000000000000000000000110100111100011111111111111111111110001111011111111111111111111110100111111110000000000000000000111001011100111111111111111111111000011101001111111111111111111100110100100010000000000000000000100101100110100000000000000000000000111110011000000000000000000010100101110101111111111111111111000100110010111111111111111111110010000011001000000000000000000010100100001010000000000000000000010001100110100000000000000000001000000100101111111111111111111101011001101000000000000000000000111101111100011111111111111111111000001111100111111111111111111110110110110100000000000000000000011111110100011111111111111111111000011011101111111111111111111111000001111000000000000000000000101111100100011111111111111111111001101010110000000000000000000001110110010011111111111111111111001111011111000000000000000000000101100010100000000000000000000010000111000010000000000000000000101001011100111111111111111111110000110100110111111111111111111101000010101001111111111111111111001001110000111111111111111111110001010011100111111111111111111111111110110111111111111111111111010010101111111111111111111111110100000010101000000000000000000011101101110001111111111111111111100001110010011111111111111111111110000000110111111111111111111111010110100000000000000000000000100101101001000000000000000000001101111100100000000000000000000010011110111101111111111111111111001010011011000000000000000000001011010111110111111111111111111100110100000111111111111111111111111001110110011111111111111111111101001100001111111111111111111101001010100001111111111111111111010111011001000000000000000000000101100110100111111111111111111111110001011111111111111111111111011000001001111111111111111111110011010011100000000000000000000011100110001101111111111111111111010010010101011111111111111111111010011010100111111111111111111101101100110101111111111111111111011100100101000000000000000000001010011111111111111111111111111100100011110110000000000000000000001010000100111111111111111111110101100110010000000000000000000000101111001011111111111111111111001001100010011111111111111111110110011101010111111111111111111100100000010010000000000000000000001101001010111111111111111111110010111001000111111111111111111111110001011110000000000000000000111111111111111111111111111111111101100100100000000000000000000001101001011010000000000000000000100011010110011111111111111111110000001011000000000000000000000000001011110100000000000000000000001110011110011111111111111111110111111011011111111111111111111100001001110001111111111111111111111101110111111111111111111111111000000011111111111111111111111101101000100001111111111111111111010000100101011111111111111111111100101010100000000000000000000001100001110011111111111111111111010001000011000000000000000000000111100100101000000000000000000011001101111001111111111111111111100100001001000000000000000000000110010011100111111111111111111100001100100000000000000000000000110010000001100000000000000000001000111001011000000000000000000001100111101010000000000000000000011111101100100000000000000000000000011000000000000000000000000001010101001101111111111111111111000011011000111111111111111111111100011111110111111111111111111111010101100000000000000000000000110110110011100000000000000000001001010100100000000000000000000000010101100111111111111111111111101011111101111111111111111111111010001110100000000000000000000011001000111011111111111111111111000010001010011111111111111111110000100111100111111111111111111110011100111000000000000000000000011001111101000000000000000000000100100000001111111111111111111110010001100000000000000000000000001111111100111111111111111111110101110011101111111111111111111110011001000000000000000000000000111011111100011111111111111111110000111000111000000000000000000011101100000001111111111111111111010000101110111111111111111111111000101001101111111111111111111100010011101111111111111111111111110010100100011111111111111111110011101110101111111111111111111101000110001111111111111111111111001100101101100000000000000000001011011011010;
    wire [32*32-1:0] bias2 = 'b1111111111111111111111101111001000000000000000000001000010100000000000000000000000001001110111010000000000000000000001101100000000000000000000000000010100010101111111111111111111111111111101010000000000000000000001110101001111111111111111111111011010101001111111111111111111011111100011111111111111111111111001110100101000000000000000000000111110001001000000000000000000001110101000000000000000000000000100011101001111111111111111111110010100000100000000000000000000001010100001100000000000000000000001000001000111111111111111111111010010010110000000000000000000001100000110111111111111111111111000001111000111111111111111111110011111111000111111111111111111100100000011110000000000000000000010110100111111111111111111111110111111111001111111111111111111110110110010101111111111111111111001011000011111111111111111111110010001001111000000000000000000000001000001111111111111111111111000000000111000000000000000000010100001000011111111111111111111110000111001001111111111111111111110001011100100000000000000000001011111011010;
    wire [32*32*16-1:0] weights3 = 'b1111111111111111111111111000101100000000000000000001000001011111000000000000000000001010010110001111111111111111110100100010100000000000000000000001101000000010000000000000000000010000010010010000000000000000001000001110011011111111111111111110010011101101111111111111111111100000110111000000000000000000001011000101100111111111111111111101111001100101000000000000000000010100100000000000000000000000000100011111001011111111111111111111100011010000111111111111111111110101110000010000000000000000001101110111010011111111111111111110101000111010111111111111111111100101001000000000000000000000001000001110110000000000000000000111111100111111000000000000000000011001110000001111111111111111111010000101111100000000000000000101011010111110000000000000000000100111001100111111111111111111111101111101101000000000000000000000010010101000000000000000000000100100011101000000000000000000001010010000000100000000000000000001101100111110000000000000000001010110100011110000000000000000000111111011100111111111111111111110001011100111111111111111111111101001010100000000000000000000000001000001001000000000000000000100000110110111000000000000000000000100001110001111111111111111111100111010111000000000000000000000011000100011000000000000000000010100011011011111111111111111111100001110111111111111111111111110101000001000111111111111111111110011010000101111111111111111110110110101111000000000000000000000101001110001000000000000000000001011011101010000000000000000000000110101010011111111111111111110010100100000000000000000000001111010001100110000000000000000001000100000110000000000000000000010001000100100000000000000000000011000101010000000000000000000100100110001001111111111111111111110110010010101000000000000000000011010010111100000000000000000110100001000010000000000000000000010100001000011111111111111111111111011000000011111111111111111111100010001100011111111111111111110010011010101111111111111111111101110111101000000000000000000010011110010000000000000000000000011110100011010000000000000000000001100001111001111111111111111110101000011101000000000000000000000011101111111111111111111111111101000001001111111111111111111101111101111000000000000000000000001001110101000000000000000000000010101011011100000000000000000000000111010010000000000000000000011000111011100111111111111111111110111101101000000000000000000000111111110011000000000000000000000100100000001000000000000000000100101111100000000000000000000000110100000000011111111111111111110111011001111111111111111111111011010100101000000000000000000000110101000000111111111111111111101101101001000111111111111111111111100010110000000000000000000001001101111101100000000000000000000000010000101111111111111111110001100001000111111111111111111111011111101010000000000000000000010011110000001111111111111111110010110110000001111111111111111111100101010001111111111111111111101100111010000111111111111111111101000001111011111111111111111111010111101000100000000000000000001001100110000111111111111111111111000101001101111111111111111100000100001001000000000000000000000110100111100111111111111111111011101010101110000000000000000001000001010110000000000000000000010000000100001111111111111111111011101000100010000000000000000000101101011100011111111111111111110100101000000111111111111111111011010000000100000000000000000000000000100011000000000000000000000000011010101111111111111111111010100101100001111111111111111111001110111111100000000000000000001110010001010000000000000000000100010101001111111111111111111111000111101011000000000000000000010001000010101111111111111111111010100111001001111111111111111111010010110101111111111111111111111000100011111000000000000000000001101011111000000000000000000001001110001011011111111111111111111110010000001111111111111111111110011111101011111111111111111111001110010001011111111111111111101111001111000000000000000000000101010101000110000000000000000000111110110010000000000000000000000100001000111111111111111111111110110110010011111111111111111111010101101111011111111111111111111101011111111000000000000000000011101101001000000000000000000000001000011011000000000000000000001010011010010000000000000000000000011100100101111111111111111111000001111011100000000000000000010100010001010000000000000000000010100111000111111111111111111111001010000000011111111111111111110011011011111111111111111111111100101010111111111111111111111111110111101101111111111111111111101111011011000000000000000000000000110110101000000000000000000001011000010100100000000000000000001100011000011000000000000000000000010110010100000000000000000000110000001010011111111111111111111001000101000111111111111111111100100101011001111111111111111111010010100011011111111111111111110001100110011111111111111111111011001011111110000000000000000001000010001101011111111111111111110110011000000000000000000000000000010010001011111111111111111111101111000101100000000000000000000011000000010111111111111111111111101100110011111111111111111111010011011010111111111111111111110001011011111111111111111111111110010010101011111111111111111110101110000010100000000000000000001010100100010000000000000000000100110000011001111111111111111110101011110101111111111111111111101100010010001000000000000000000010011100001100000000000000000000000001101011111111111111111111111111110001110000000000000000000100101111001011111111111111111111010011001101100000000000000000010010100011011111111111111111111011011101111010000000000000000000101110000010000000000000000000000111100001110111111111111111111100001010101111111111111111111111010010101101100000000000000000001001010011101111111111111111111010110101000111111111111111111111001110001011011111111111111111101010100100011111111111111111111111110110011100000000000000000000001111100110011111111111111111101110101000111000000000000000000100100100100111111111111111111111010101001011011111111111111111101111010001111111111111111111111100000000010100000000000000000000111101110000100000000000000000001111010010001000000000000000000011000000101111111111111111111111111101110101000000000000000000000000101111101000000000000000000011000110110011111111111111111111010001010001011111111111111111111000001110001000000000000000000011111110100011111111111111111111000111010011111111111111111111101101000100010111111111111111111110011001110010000000000000000001000101000000111111111111111111111110111011001000000000000000000000011010100111111111111111111110101011111000000000000000000000000110111100101111111111111111111100001011011011111111111111111111100100111001100000000000000000001000110111010111111111111111111100010011010010000000000000000001010010100010100000000000000000000001000011000111111111111111111100011011000011111111111111111111110001001000100000000000000000001111011011100111111111111111111111100110101110000000000000000001010110100100100000000000000000010100111010111000000000000000000011001111111011111111111111111111000001011000111111111111111111101100101011000000000000000000000100010101000001111111111111111110110001100011111111111111111111111001010001111111111111111111111101111011010110000000000000000000110000110110100000000000000000010010011001001111111111111111111110001011010000000000000000000000010000000010111111111111111111101010000011001000000000000000000010010001100001111111111111111111100001110011111111111111111111111101111001110000000000000000000011001000000010000000000000000000100000011100011111111111111111111000111010011000000000000000000001110010110000000000000000000000001111110000100000000000000000001001011110001000000000000000000011111110100110000000000000000000010111010111100000000000000000000010100000011111111111111111111011100110010000000000000000000000010010011001011111111111111111110111111101111000000000000000000010100100110111111111111111111110110101011001111111111111111111111010110011010111111111111111111010101000000001111111111111111111010001101100011111111111111111111011101111000111111111111111111100000011100111111111111111111111100110110111100000000000000000000101111111101000000000000000000101011001110000000000000000000001000011110100111111111111111111111001010001001000000000000000000010000100000111111111111111111111000111000100111111111111111111110011110001100000000000000000000100111101011000000000000000000000110001000001100000000000000000000101001001000111111111111111111101011110001101111111111111111110101100011110111111111111111111111010111110111111111111111111111111000101010010000000000000000000001111010011000000000000000000001101011010011000000000000000000010110011001100000000000000000001010110100010111111111111111111111101100011000000000000000000000010011111111001111111111111111111011110000101011111111111111111111001110011001111111111111111111100010011100001111111111111111110110111101110111111111111111111101001010111100111111111111111111110011101101001111111111111111111011011100100100000000000000000010100100000110000000000000000000101001110111100000000000000000000101001001011011111111111111111110011011111001111111111111111111011001011101001111111111111111111011110101001011111111111111111111100111101100111111111111111111110011011101100000000000000000000101010011100000000000000000000001010010101001111111111111111111010101111010001111111111111111101111110110000100000000000000000000100111111100000000000000000000011011101101000000000000000000001101101000001111111111111111111110101010110110000000000000000000100111110111011111111111111111110101111100101011111111111111111111000110110001111111111111111111110111110001011111111111111111110101001100001111111111111111111111010001100110111111111111111111110001010010100000000000000000000110000000111100000000000000000001000101001000000000000000000000010111011110100000000000000000000110010000010111111111111111111111001010011100111111111111111111100111010110010000000000000000011000101000100000000000000000000010101101010010000000000000000000011100001101011111111111111111110101101110100100000000000000001000100001011010000000000000000000101100010011011111111111111111111110000100000100000000000000000101111100010001000000000000000000100011010011011111111111111111110101000011110100000000000000000001100110100101111111111111111111110001001011100000000000000000000011010100011000000000000000000100110101000011000000000000000001000110000101000000000000000000001010100011100100000000000000000001101110100000000000000000000000010011000001110000000000000000000111011110011011111111111111111101010000111000111111111111111111100000101011100000000000000000000010001000100111111111111111111111010110011111111111111111111111110101111101101111111111111111111011001001011000000000000000000010100101101001111111111111111111100011100111010000000000000000000100110110101000000000000000000000001011100100000000000000000000001010001001111111111111111111110101111110001011111111111111111110010011010000000000000000000000000100111111101111111111111111111011000110000100000000000000000000100000010101000000000000000000100100011000110000000000000000000000001111000011111111111111111110111001010101111111111111111111110000110010010000000000000000000001100101000011111111111111111101110000110111000000000000000000010010000010010000000000000000001001101100001111111111111111111101111100100110000000000000000000000101100001010000000000000000001000011110000000000000000000000001101001001100000000000000000000001001110000111111111111111111110101111111001000000000000000000000011110101000111111111111111111110001110000110000000000000000000000011000101111111111111111111110001010010000111111111111111111011110001101000000000000000000000001001011000011111111111111111101010011001110111111111111111111011010100010110000000000000000001010111000101011111111111111111101101011001101111111111111111111011110100100001111111111111111110011010111101111111111111111111110010101111011000000000000000000011011001110010000000000000000000101000100000111111111111111111110000011101011111111111111111111100100010011110000000000000000001001001001001111111111111111111101110000000110111111111111111111011010001011001111111111111111111001000000001100000000000000000010001101111111000000000000000000011101011110011111111111111111111111110111000011111111111111111111000011100110000000000000000000001010011110011111111111111111110100101100001011111111111111111101111001010101000000000000000000010011111010010000000000000000000111011110100000000000000000000001010111001010000000000000000000101001110011001111111111111111101110110111111000000000000000000000110000010101000000000000000000101010010001101111111111111111111000111001001100000000000000000010101101111010111111111111111111111000001101100000000000000000000000010111111100000000000000000001110001100000000000000000000000011010000111111111111111111111111100001001111100000000000000000000101001110101111111111111111111011011100111110000000000000000001011000111101000000000000000000010000111000010111111111111111111110111011011000000000000000000000111001001110011111111111111111101111000110010111111111111111111100101001010100000000000000000001001100100101111111111111111111011110101010111000000000000000000000110011111000000000000000000000000010110101100000000000000000001010000010010111111111111111111000010101010010000000000000000000100100101101100000000000000000000011000101101111111111111111111110100100011000000000000000000000001101010011011111111111111111100100000111000000000000000000000100010110010001111111111111111111011110111110100000000000000000001111010000111111111111111111111011101101010001111111111111111111111110110010011111111111111111110101010100010111111111111111111110000111011100000000000000000000011001010100000000000000000000000111000101110000000000000000000001111011100000000000000000000000000010001111000000000000000000000011001101110111111111111111111111010001001000000000000000000001001010001000111111111111111111101110101011111111111111111111111110111001111110000000000000000000000110000000000000000000000000000001110010010000000000000000000010111010100001111111111111111111101101011011011111111111111111101001111010000111111111111111111011100000001001111111111111111111011000111011111111111111111111100111100000110111111111111111111100110001010001111111111111111111011011100001111111111111111111110010010000000111111111111111111010110000100101111111111111111111100111100101011111111111111111101111101001100111111111111111111110000101001101111111111111111111110100100001000000000000000000000010110010001111111111111111111111011001110110000000000000000000110010001011000000000000000000001100100111011000000000000000000001000111111010000000000000000001011010111111000000000000000000001111001010100000000000000000000000000001101000000000000000000000000000101011011111111111111111101110011110101111111111111111111100110101111001111111111111111111100010111011100000000000000000010101010011011111111111111111111111001110011010000000000000000000101010100011011111111111111111111101011000101000000000000000000101101010111001111111111111111111110101000010100000000000000000101011011010010111111111111111111110100000101100000000000000000000101010110011011111111111111111110010101101000000000000000000001011010100001100000000000000000000011111101011011111111111111111101111100111011000000000000000001001010101100010000000000000000001100001111011011111111111111111111101101001101000000000000000000101010010111110000000000000000001000111111100011111111111111111111001011001011000000000000000000111010111110110000000000000000011010000110110111111111111111111110010010000000111111111111111111111011110100010000000000000000001101010010110011111111111111111110000100010010000000000000000000010001111100110000000000000000001001110111010011111111111111111111101110000001000000000000000000101110000000110000000000000000000000001010110000000000000000000000100011101111111111111111111111101111100001101111111111111111111011001100001000000000000000000010001001100001000000000000000000010010000010011111111111111111111110010100111111111111111111111111100111110011000000000000000000000011000000001111111111111111110111001010010111111111111111111110111110100110000000000000000000001001110001100000000000000000001000111010111100000000000000000001000110010110111111111111111111011111100001011111111111111111110011111100011011111111111111111111111000001100000000000000000000101100000111111111111111111111111110001101111100000000000000000000111011100101111111111111111111110001001101010000000000000000001010111000110000000000000000000011010000010110000000000000000000010101001101100000000000000000000111100100000000000000000000000000000110010101;
    wire [32*16-1:0] bias3 = 'b11111111111111111111101010011111111111111111111111101101110010000000000000000000001001111000010000000000000000000010110100111111111111111111111111011111010001001111111111111111110111110001101000000000000000000000000000010011111111111111111111101010000010001111111111111111111101110101110111111111111111111111111111001000000000000000000000000100100101001111111111111111111001101110101100000000000000000001110110011001000000000000000000010100101010000000000000000000000101000000010100000000000000000000001100111000;
    wire [32*16-1:0] weights4 ='b00000000000000000010111010001100000000000000000001000100001011101111111111111111110100110100011011111111111111111111110010111100111111111111111111011010000100101111111111111111111100000010110100000000000000000010111111000110000000000000000000011010001001100000000000000000000110001110101000000000000000000101110100000001111111111111111111001010001001011111111111111111110100111011111111111111111111111100001011000001111111111111111111111010110110110000000000000000010011000100010111111111111111111001011100110001;
    wire [32-1:0] bias4 = 'b11111111111111111111010010100111;

    //testing inputs
    //entry 75 of spreadsheet
    //wire [127:0] in_data1 = 'b00000000000000101100000000011010000000111110011011001100110011010000010010110010110101011000100000001011101111111011111000001111; 
    //entry 12 
    //wire [127:0] in_data1 = 'b00000000000000100110010100101100000000111110011100000000000000000000000010100110011110111101101000000001100011001010001100110011; 
    //entry 64
    wire [127:0] in_data1 = 'b00000000000000101001111111010010000000111110011011001100110011010000010000001000001011111111100100001001111110010001110111010011;  
    //entry 97588
    //wire [127:0] in_data1 = 'b00000000000000101100000000000111000000111110011011001100110011010000001001100110011000000101010000000110000111000111000111100110;  
    
	// Instantiate the prediction module
    battery_soh_predictor predictor (
        .clk(clk),
        .reset(reset),
        .in_data(in_data1),
        .weights1(weights1),
        .bias1(bias1),
        .weights2(weights2),
        .bias2(bias2),
        .weights3(weights3),
        .bias3(bias3),
        .weights4(weights4),
        .bias4(bias4),
        .soh_out(predicted_soh)
    );
    
endmodule
